`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:			
//					
// Engineer: 		
//
// Create Date:		
// Design Name: 	
// Module Name:     
// Project Name:	
// Target Devices: 
// Tool versions:
// Description:		
//
// Dependencies:
//
// Revision:
//
//
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module program_counter
(
    //--------------------------
	// Input Ports
	//--------------------------
	input				clk,
	input				rst,
	input		[3:0]	pc_control,
	input		[25:0]	jump_address,
	input		[15:0]	branch_offset,
	input		[31:0] 	reg_address,
	
    //--------------------------
    // Output Ports
    //--------------------------
    output 	reg	[31:0] 	pc

); 
      
    ///////////////////////////////////////////////////////////////////
    // Begin Design
    ///////////////////////////////////////////////////////////////////
    //-------------------------------------------------
    // Signal Declarations: local params
    //-------------------------------------------------
   
    //-------------------------------------------------
    // Signal Declarations: reg
    //-------------------------------------------------    
	
    //-------------------------------------------------
    // Signal Declarations: wire
    //-------------------------------------------------
	
	//---------------------------------------------------------------
	// Instantiations
	//---------------------------------------------------------------
	// None

	//---------------------------------------------------------------
	// Combinatorial Logic
	//---------------------------------------------------------------
		
	//---------------------------------------------------------------
	// Sequential Logic
	//---------------------------------------------------------------
	
	always @(posedge clk or posedge rst)
	begin
		if (rst)
		begin
			pc <= 32'd0;
		end
		else
		begin
			case (pc_control)
				4'b0000 : pc <= pc + 32'd4;
				4'b0001 : pc <= {pc[31:28],(jump_address[25:0]),2'b00};
				4'b0010 : pc <= reg_address;
				4'b0011 : pc <= pc + 32'd4 + ({{16{branch_offset[15]}},branch_offset} << 2);
				default : pc <= pc;
			endcase
		end
	end
    
 endmodule  



