`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:			
//					
// Engineer: 		
//
// Create Date:		
// Design Name: 	
// Module Name:     
// Project Name:	
// Target Devices: 
// Tool versions:
// Description:		
//
// Dependencies:
//
// Revision:
//
//
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module mux_2to1

(
    in0,	//input 0
	in1,	//input 1
	out,	//output
	sel	//select
);

    //--------------------------
	// Parameters
	//--------------------------	
	parameter DWIDTH = 32;
    //--------------------------
	// Input Ports
	//--------------------------
	// < Enter Input Ports  >
    input 		[DWIDTH-1:0]		in0;
	input 		[DWIDTH-1:0]		in1;
	input 									sel;
	
    //--------------------------
    // Output Ports
    //--------------------------
    // < Enter Output Ports  >	
    output 	[DWIDTH-1:0] 		out; 
		
    //--------------------------
    // Bidirectional Ports
    //--------------------------
    // < Enter Bidirectional Ports in Alphabetical Order >
    // None
      
    ///////////////////////////////////////////////////////////////////
    // Begin Design
    ///////////////////////////////////////////////////////////////////
    //-------------------------------------------------
    // Signal Declarations: local params
    //-------------------------------------------------
   
    //-------------------------------------------------
    // Signal Declarations: reg
    //-------------------------------------------------    
    
    //-------------------------------------------------
    // Signal Declarations: wire
    //-------------------------------------------------
		
	//---------------------------------------------------------------
	// Instantiations
	//---------------------------------------------------------------
	// None

	//---------------------------------------------------------------
	// Combinatorial Logic
	//---------------------------------------------------------------
	assign out = (sel == 0) ? in0 : in1;
	
	//---------------------------------------------------------------
	// Sequential Logic
	//---------------------------------------------------------------
    
 endmodule  



